// 2022.09.05

module Q10172();
    initial begin
        $display("|\\_/|");
        $display("|q p|   /}");
        $display("( 0 )\"\"\"\\");
        $display("|\"^\"`    |");
        $display("||_/=\\\\__|");
        $finish;
    end
endmodule