// 2022.09.05

module Q10171();
    initial begin
        $display("\\    /\\");
        $display(" )  ( ')");
        $display("(  /  )");
        $display(" \\(__)|");
        $finish;
    end
endmodule