// 2022.09.05

module Q25083();
    initial begin
        $display("         ,r'\"7");
        $display("r`-_   ,'  ,/");
        $display(" \\. \". L_r'");
        $display("   `~\\/");
        $display("      |");
        $display("      |");
        $finish;
    end
endmodule