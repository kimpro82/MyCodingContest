// 2022.08.18

module Q2557();
    initial begin
        $display("Hello World!");
        $finish;
    end
endmodule