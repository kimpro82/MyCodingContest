// 2022.09.05

module Q10718();

    initial begin
        repeat (2) begin
            $display("강한친구 대한육군");
        end
        $finish;
    end

endmodule